module MAIN_DECODER 
(
    input wire [4:0] Opcode,
    output red       MemtoReg,
    output red       MemWrite,
    output red       Branch,
    output red       ALUSrc,
);
    
endmodule